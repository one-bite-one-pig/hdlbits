module top_module(
    input clk,
    input areset,    // Freshly brainwashed Lemmings walk left.
    input bump_left,
    input bump_right,
    output walk_left,
    output walk_right); //  

    parameter LEFT=0, RIGHT=1;
    reg state, next_state;

    always @(*) begin
        // State transition logic
        if (state==0)begin
            if(bump_left) next_state=RIGHT;
            else next_state=LEFT;
        end
        else begin
            if(bump_right) next_state=LEFT;
            else next_state=RIGHT;
        end
    end

    always @(posedge clk, posedge areset) begin
        // State flip-flops with asynchronous reset
        if(areset) state<=LEFT;
        else state<=next_state;
    end

    
    assign walk_left = (state == LEFT);
    assign walk_right = (state == RIGHT);

endmodule