module top_module(
    input [31:0] a,
    input [31:0] b,
    output [31:0] sum
);
    wire c1;
    wire[16:0] h1,h2;
    add16 m1(.a(a[15:0]),.b(b[15:0]),.cin(1'b0),.cout(c1),.sum(sum[15:0]));
    add16 m2(.a(a[31:16]),.b(b[31:16]),.cin(1'b0),.sum(h1));
    add16 m3(.a(a[31:16]),.b(b[31:16]),.cin(1'b1),.sum(h2));
    assign sum[31:16]=c1? h2:h1;

endmodule